module systolic_mult(); 

    input 